module top_module(
    input a, 
    input b,
    output wire out_assign,
    output reg out_alwaysblock
);

endmodule